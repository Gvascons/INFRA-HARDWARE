module StoreBlock(
	input logic [63:0]Entrada,
	input logic [2:0]StoreTYPE,
	output logic [63:0]StoreResult);
	
	always_comb begin
	
	end
endmodule //LoadBlock





